`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Cal Poly SLO CPE 133
// Engineer: Darian Primer
// 
// Create Date: 10/11/2018 10:35:08 AM 
// Description: Lab 3 SIM file
//////////////////////////////////////////////////////////////////////////////////


module Lab3SIM();

logic [3:0] A, B;
logic [3:0] an;
logic [6:0] sseg;

Lab3 Lab3_inst(.*);




endmodule
